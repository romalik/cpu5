// Hex inverter

module ttl_7404 #(parameter BLOCKS = 6, DELAY_RISE = 0, DELAY_FALL = 0)
(
  input [BLOCKS-1:0] A,
  output [BLOCKS-1:0] Y
);
/*verilator inline_module*/
//------------------------------------------------//
reg [BLOCKS-1:0] computed;

always @(*)
begin
  computed = ~A;
end
//------------------------------------------------//

assign Y = computed;

endmodule
